typedef struct {
  logic[31:0] a;
  logic[31:0] b;
  logic[31:0] c;
  logic[31:0] d;
  logic[31:0] e;
  logic[31:0] f;
  logic[31:0] g;
  logic[31:0] h;
} HashState;
