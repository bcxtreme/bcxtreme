
module golden_sha_stim();

  golden_sha test;

endmodule

